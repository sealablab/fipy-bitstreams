library IEEE;
use IEEE.Std_Logic_1164.all;
use IEEE.Numeric_Std.all;


architecture Behavioural of CustomWrapper is
begin
    -- ___ <= InputA;
    -- ___ <= InputB;
    -- ___ <= InputC;
    -- ___ <= InputD;

    -- ___ <= Control0;
    -- ___ <= Control1;
    -- ___ <= Control2;
    --      ...
    -- ___ <= Control15;

    -- OutputA => ___;
    -- OutputB => ___;
    -- OutputC => ___;
    -- OutputD => ___;
end architecture;
