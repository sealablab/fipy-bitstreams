library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rom_slow is
    generic (
        rom_width: integer := 10
    );
	Port (
		clk : in STD_LOGIC;
		address : in STD_LOGIC_VECTOR(15 downto 0);
		data_out : out STD_LOGIC_VECTOR(15 downto 0)
	);
end rom_slow;

architecture Behavioral of rom_slow is

type romtype is array(0 to 2**rom_width-1) of std_logic_vector(15 downto 0);    

  signal memory_ram : romtype := (x"0001", x"0002", x"0003", x"0004", x"0005", x"0006", x"0007", x"0008", x"0009", x"000a", x"000b", x"000c", x"000d", x"000e", x"000f", x"0010", x"0011", x"0012", x"0013", x"0014", x"0015", x"0016", x"0017", x"0018", x"0019", x"001a", x"001b", x"001c", x"001d", x"001e", x"001f", x"0020", x"0021", x"0022", x"0023", x"0024", x"0025", x"0026", x"0027", x"0028", x"0029", x"002a", x"002b", x"002c", x"002d", x"002e", x"002f", x"0030", x"0031", x"0032", x"0033", x"0034", x"0035", x"0036", x"0037", x"0038", x"0039", x"003a", x"003b", x"003c", x"003d", x"003e", x"003f", x"0040", x"0041", x"0042", x"0043", x"0044", x"0045", x"0046", x"0047", x"0048", x"0049", x"004a", x"004b", x"004c", x"004d", x"004e", x"004f", x"0050", x"0051", x"0052", x"0053", x"0054", x"0055", x"0056", x"0057", x"0058", x"0059", x"005a", x"005b", x"005c", x"005d", x"005e", x"005f", x"0060", x"0061", x"0062", x"0063", x"0064", x"0065", x"0066", x"0067", x"0068", x"0069", x"006a", x"006b", x"006c", x"006d", x"006e", x"006f", x"0070", x"0071", x"0072", x"0073", x"0074", x"0075", x"0076", x"0077", x"0078", x"0079", x"007a", x"007b", x"007c", x"007d", x"007e", x"007f", 
x"0080", x"0081", x"0082", x"0083", x"0084", x"0085", x"0086", x"0087", x"0088", x"0089", x"008a", x"008b", x"008c", x"008d", x"008e", x"008f", x"0090", x"0091", x"0092", x"0093", x"0094", x"0095", x"0096", x"0097", x"0098", x"0099", x"009a", x"009b", x"009c", x"009d", x"009e", x"009f", x"00a0", x"00a1", x"00a2", x"00a3", x"00a4", x"00a5", x"00a6", x"00a7", x"00a8", x"00a9", x"00aa", x"00ab", x"00ac", x"00ad", x"00ae", x"00af", x"00b0", x"00b1", x"00b2", x"00b3", x"00b4", x"00b5", x"00b6", x"00b7", x"00b8", x"00b9", x"00ba", x"00bb", x"00bc", x"00bd", x"00be", x"00bf", x"00c0", x"00c1", x"00c2", x"00c3", x"00c4", x"00c5", x"00c6", x"00c7", x"00c8", x"00c9", x"00ca", x"00cb", x"00cc", x"00cd", x"00ce", x"00cf", x"00d0", x"00d1", x"00d2", x"00d3", x"00d4", x"00d5", x"00d6", x"00d7", x"00d8", x"00d9", x"00da", x"00db", x"00dc", x"00dd", x"00de", x"00df", x"00e0", x"00e1", x"00e2", x"00e3", x"00e4", x"00e5", x"00e6", x"00e7", x"00e8", x"00e9", x"00ea", x"00eb", x"00ec", x"00ed", x"00ee", x"00ef", x"00f0", x"00f1", x"00f2", x"00f3", x"00f4", x"00f5", x"00f6", x"00f7", x"00f8", x"00f9", x"00fa", x"00fb", x"00fc", x"00fd", x"00fe", x"00ff", 
x"0100", x"0101", x"0102", x"0103", x"0104", x"0105", x"0106", x"0107", x"0108", x"0109", x"010a", x"010b", x"010c", x"010d", x"010e", x"010f", x"0110", x"0111", x"0112", x"0113", x"0114", x"0115", x"0116", x"0117", x"0118", x"0119", x"011a", x"011b", x"011c", x"011d", x"011e", x"011f", x"0120", x"0121", x"0122", x"0123", x"0124", x"0125", x"0126", x"0127", x"0128", x"0129", x"012a", x"012b", x"012c", x"012d", x"012e", x"012f", x"0130", x"0131", x"0132", x"0133", x"0134", x"0135", x"0136", x"0137", x"0138", x"0139", x"013a", x"013b", x"013c", x"013d", x"013e", x"013f", x"0140", x"0141", x"0142", x"0143", x"0144", x"0145", x"0146", x"0147", x"0148", x"0149", x"014a", x"014b", x"014c", x"014d", x"014e", x"014f", x"0150", x"0151", x"0152", x"0153", x"0154", x"0155", x"0156", x"0157", x"0158", x"0159", x"015a", x"015b", x"015c", x"015d", x"015e", x"015f", x"0160", x"0161", x"0162", x"0163", x"0164", x"0165", x"0166", x"0167", x"0168", x"0169", x"016a", x"016b", x"016c", x"016d", x"016e", x"016f", x"0170", x"0171", x"0172", x"0173", x"0174", x"0175", x"0176", x"0177", x"0178", x"0179", x"017a", x"017b", x"017c", x"017d", x"017e", x"017f", 
x"0180", x"0181", x"0182", x"0183", x"0184", x"0185", x"0186", x"0187", x"0188", x"0189", x"018a", x"018b", x"018c", x"018d", x"018e", x"018f", x"0190", x"0191", x"0192", x"0193", x"0194", x"0195", x"0196", x"0197", x"0198", x"0199", x"019a", x"019b", x"019c", x"019d", x"019e", x"019f", x"01a0", x"01a1", x"01a2", x"01a3", x"01a4", x"01a5", x"01a6", x"01a7", x"01a8", x"01a9", x"01aa", x"01ab", x"01ac", x"01ad", x"01ae", x"01af", x"01b0", x"01b1", x"01b2", x"01b3", x"01b4", x"01b5", x"01b6", x"01b7", x"01b8", x"01b9", x"01ba", x"01bb", x"01bc", x"01bd", x"01be", x"01bf", x"01c0", x"01c1", x"01c2", x"01c3", x"01c4", x"01c5", x"01c6", x"01c7", x"01c8", x"01c9", x"01ca", x"01cb", x"01cc", x"01cd", x"01ce", x"01cf", x"01d0", x"01d1", x"01d2", x"01d3", x"01d4", x"01d5", x"01d6", x"01d7", x"01d8", x"01d9", x"01da", x"01db", x"01dc", x"01dd", x"01de", x"01df", x"01e0", x"01e1", x"01e2", x"01e3", x"01e4", x"01e5", x"01e6", x"01e7", x"01e8", x"01e9", x"01ea", x"01eb", x"01ec", x"01ed", x"01ee", x"01ef", x"01f0", x"01f1", x"01f2", x"01f3", x"01f4", x"01f5", x"01f6", x"01f7", x"01f8", x"01f9", x"01fa", x"01fb", x"01fc", x"01fd", x"01fe", x"01ff", 
x"0200", x"0201", x"0202", x"0203", x"0204", x"0205", x"0206", x"0207", x"0208", x"0209", x"020a", x"020b", x"020c", x"020d", x"020e", x"020f", x"0210", x"0211", x"0212", x"0213", x"0214", x"0215", x"0216", x"0217", x"0218", x"0219", x"021a", x"021b", x"021c", x"021d", x"021e", x"021f", x"0220", x"0221", x"0222", x"0223", x"0224", x"0225", x"0226", x"0227", x"0228", x"0229", x"022a", x"022b", x"022c", x"022d", x"022e", x"022f", x"0230", x"0231", x"0232", x"0233", x"0234", x"0235", x"0236", x"0237", x"0238", x"0239", x"023a", x"023b", x"023c", x"023d", x"023e", x"023f", x"0240", x"0241", x"0242", x"0243", x"0244", x"0245", x"0246", x"0247", x"0248", x"0249", x"024a", x"024b", x"024c", x"024d", x"024e", x"024f", x"0250", x"0251", x"0252", x"0253", x"0254", x"0255", x"0256", x"0257", x"0258", x"0259", x"025a", x"025b", x"025c", x"025d", x"025e", x"025f", x"0260", x"0261", x"0262", x"0263", x"0264", x"0265", x"0266", x"0267", x"0268", x"0269", x"026a", x"026b", x"026c", x"026d", x"026e", x"026f", x"0270", x"0271", x"0272", x"0273", x"0274", x"0275", x"0276", x"0277", x"0278", x"0279", x"027a", x"027b", x"027c", x"027d", x"027e", x"027f", 
x"0280", x"0281", x"0282", x"0283", x"0284", x"0285", x"0286", x"0287", x"0288", x"0289", x"028a", x"028b", x"028c", x"028d", x"028e", x"028f", x"0290", x"0291", x"0292", x"0293", x"0294", x"0295", x"0296", x"0297", x"0298", x"0299", x"029a", x"029b", x"029c", x"029d", x"029e", x"029f", x"02a0", x"02a1", x"02a2", x"02a3", x"02a4", x"02a5", x"02a6", x"02a7", x"02a8", x"02a9", x"02aa", x"02ab", x"02ac", x"02ad", x"02ae", x"02af", x"02b0", x"02b1", x"02b2", x"02b3", x"02b4", x"02b5", x"02b6", x"02b7", x"02b8", x"02b9", x"02ba", x"02bb", x"02bc", x"02bd", x"02be", x"02bf", x"02c0", x"02c1", x"02c2", x"02c3", x"02c4", x"02c5", x"02c6", x"02c7", x"02c8", x"02c9", x"02ca", x"02cb", x"02cc", x"02cd", x"02ce", x"02cf", x"02d0", x"02d1", x"02d2", x"02d3", x"02d4", x"02d5", x"02d6", x"02d7", x"02d8", x"02d9", x"02da", x"02db", x"02dc", x"02dd", x"02de", x"02df", x"02e0", x"02e1", x"02e2", x"02e3", x"02e4", x"02e5", x"02e6", x"02e7", x"02e8", x"02e9", x"02ea", x"02eb", x"02ec", x"02ed", x"02ee", x"02ef", x"02f0", x"02f1", x"02f2", x"02f3", x"02f4", x"02f5", x"02f6", x"02f7", x"02f8", x"02f9", x"02fa", x"02fb", x"02fc", x"02fd", x"02fe", x"02ff", 
x"0300", x"0301", x"0302", x"0303", x"0304", x"0305", x"0306", x"0307", x"0308", x"0309", x"030a", x"030b", x"030c", x"030d", x"030e", x"030f", x"0310", x"0311", x"0312", x"0313", x"0314", x"0315", x"0316", x"0317", x"0318", x"0319", x"031a", x"031b", x"031c", x"031d", x"031e", x"031f", x"0320", x"0321", x"0322", x"0323", x"0324", x"0325", x"0326", x"0327", x"0328", x"0329", x"032a", x"032b", x"032c", x"032d", x"032e", x"032f", x"0330", x"0331", x"0332", x"0333", x"0334", x"0335", x"0336", x"0337", x"0338", x"0339", x"033a", x"033b", x"033c", x"033d", x"033e", x"033f", x"0340", x"0341", x"0342", x"0343", x"0344", x"0345", x"0346", x"0347", x"0348", x"0349", x"034a", x"034b", x"034c", x"034d", x"034e", x"034f", x"0350", x"0351", x"0352", x"0353", x"0354", x"0355", x"0356", x"0357", x"0358", x"0359", x"035a", x"035b", x"035c", x"035d", x"035e", x"035f", x"0360", x"0361", x"0362", x"0363", x"0364", x"0365", x"0366", x"0367", x"0368", x"0369", x"036a", x"036b", x"036c", x"036d", x"036e", x"036f", x"0370", x"0371", x"0372", x"0373", x"0374", x"0375", x"0376", x"0377", x"0378", x"0379", x"037a", x"037b", x"037c", x"037d", x"037e", x"037f", 
x"0380", x"0381", x"0382", x"0383", x"0384", x"0385", x"0386", x"0387", x"0388", x"0389", x"038a", x"038b", x"038c", x"038d", x"038e", x"038f", x"0390", x"0391", x"0392", x"0393", x"0394", x"0395", x"0396", x"0397", x"0398", x"0399", x"039a", x"039b", x"039c", x"039d", x"039e", x"039f", x"03a0", x"03a1", x"03a2", x"03a3", x"03a4", x"03a5", x"03a6", x"03a7", x"03a8", x"03a9", x"03aa", x"03ab", x"03ac", x"03ad", x"03ae", x"03af", x"03b0", x"03b1", x"03b2", x"03b3", x"03b4", x"03b5", x"03b6", x"03b7", x"03b8", x"03b9", x"03ba", x"03bb", x"03bc", x"03bd", x"03be", x"03bf", x"03c0", x"03c1", x"03c2", x"03c3", x"03c4", x"03c5", x"03c6", x"03c7", x"03c8", x"03c9", x"03ca", x"03cb", x"03cc", x"03cd", x"03ce", x"03cf", x"03d0", x"03d1", x"03d2", x"03d3", x"03d4", x"03d5", x"03d6", x"03d7", x"03d8", x"03d9", x"03da", x"03db", x"03dc", x"03dd", x"03de", x"03df", x"03e0", x"03e1", x"03e2", x"03e3", x"03e4", x"03e5", x"03e6", x"03e7", x"03e8", x"03e9", x"03ea", x"03eb", x"03ec", x"03ed", x"03ee", x"03ef", x"03f0", x"03f1", x"03f2", x"03f3", x"03f4", x"03f5", x"03f6", x"03f7", x"03f8", x"03f9", x"03fa", x"03fb", x"03fc", x"03fd", x"03fe", x"03ff", 
x"0400");

begin                                                        

process (clk)                                                
begin                                                        
	if(rising_edge(clk)) then  
		data_out <= memory_ram(to_integer(unsigned(address)));      
	end if;                                                      
end process;             

end Behavioral;